module dut (P1, P2, P3, P4);

  input P1, P2;
  output [7:0] P3;
  inout P4;
  
endmodule