module sample(
    clk,
    rst,
    data_i,
    data_o
);

// input & output
input clk;
input rst;
input data_i;
output data_o;

endmodule
