package dummy_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "dummy_if.sv"
  `include "dummy_item.sv"
  `include "dummy_driver.sv"
  `include "dummy_monitor.sv"
  `include "dummy_agent.sv"
  `include "dummy_env.sv"

endpackage: dummy_pkg
